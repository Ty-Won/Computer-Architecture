LIBRARY ieee;
USE ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

ENTITY pipeline_tb IS
END pipeline_tb;

ARCHITECTURE behaviour OF pipeline_tb IS

COMPONENT pipeline IS
port (clk : in std_logic;
      a, b, c, d, e : in integer;
      op1, op2, op3, op4, op5, final_output : out integer
  );
END COMPONENT;

--The input signals with their initial values
SIGNAL clk: STD_LOGIC := '0';
SIGNAL s_a, s_b, s_c, s_d, s_e : INTEGER := 0;
SIGNAL s_op1, s_op2, s_op3, s_op4, s_op5, s_final_output : INTEGER := 0;

CONSTANT clk_period : time := 1 ns;

BEGIN
dut: pipeline
PORT MAP(clk, s_a, s_b, s_c, s_d, s_e, s_op1, s_op2, s_op3, s_op4, s_op5, s_final_output);

 --clock process
clk_process : PROCESS
BEGIN
	clk <= '0';
	WAIT FOR clk_period/2;
	clk <= '1';
	WAIT FOR clk_period/2;
END PROCESS;
 

stim_process: PROCESS
BEGIN   
	-- FULL
	REPORT "Filling up pipeline with full input [a=1,b=2,c=3,d=4,e=5]";
	s_a <= 1;
	s_b <= 2;
	s_c <= 3;
	s_d <= 4;
	s_e <= 5;
	WAIT FOR 1 * clk_period;
	ASSERT (s_op1 = 3) REPORT "the output should be '3'" SEVERITY ERROR;
	ASSERT (s_op2 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op3 = 12) REPORT "the output should be '12'" SEVERITY ERROR;
	ASSERT (s_op4 = -4) REPORT "the output should be '-4'" SEVERITY ERROR;
	ASSERT (s_op5 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_final_output = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	REPORT "_______________________";


	REPORT "Filling up pipeline with another input [a=5,b=2,c=4,d=10,e=6]";
	s_a <= 5;
	s_b <= 2;
	s_c <= 4;
	s_d <= 10;
	s_e <= 6;
	WAIT FOR 1 * clk_period;
	ASSERT (s_op1 = 7) REPORT "the output should be '7'" SEVERITY ERROR;
	ASSERT (s_op2 = 126) REPORT "the output should be '126'" SEVERITY ERROR;
	ASSERT (s_op3 = 40) REPORT "the output should be '40'" SEVERITY ERROR;
	ASSERT (s_op4 = -1) REPORT "the output should be '-1'" SEVERITY ERROR;
	ASSERT (s_op5 = -48) REPORT "the output should be '-48'" SEVERITY ERROR;
	ASSERT (s_final_output = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	REPORT "_______________________";


	REPORT " Filling up pipeline with another input[a=0,b=3,c=1,d=2,e=2]";
	s_a <= 0;
	s_b <= 3;
	s_c <= 1;
	s_d <= 2;
	s_e <= 2;
	WAIT FOR 1 * clk_period;
	ASSERT (s_op1 = 3) REPORT "the output should be '3'" SEVERITY ERROR;
	ASSERT (s_op2 = 294) REPORT "the output should be '294'" SEVERITY ERROR;
	ASSERT (s_op3 = 2) REPORT "the output should be '2'" SEVERITY ERROR;
	ASSERT (s_op4 = -2) REPORT "the output should be '-2'" SEVERITY ERROR;
	ASSERT (s_op5 = -40) REPORT "the output should be '-40'" SEVERITY ERROR;
	ASSERT (s_final_output = 174) REPORT "the output should be '174'" SEVERITY ERROR;
	REPORT "_______________________";

	--half full
	REPORT "Begin draining the pipeline to make it half full [a=0,b=0,c=0,d=0,e=0]";
	s_a <= 0;
	s_b <= 0;
	s_c <= 0;
	s_d <= 0;
	s_e <= 0;
	WAIT FOR 1 * clk_period;
	ASSERT (s_op1 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op2 = 126) REPORT "the output should be '126'" SEVERITY ERROR;
	ASSERT (s_op3 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op4 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op5 = -4) REPORT "the output should be '-40'" SEVERITY ERROR;
	ASSERT (s_final_output = 334) REPORT "the output should be '334'" SEVERITY ERROR;
	REPORT "_______________________";


	--emptying the pipeline
	REPORT "Draining the pipeline [a=0,b=0,c=0,d=0,e=0]";
	s_a <= 0;
	s_b <= 0;
	s_c <= 0;
	s_d <= 0;
	s_e <= 0;
	WAIT FOR 1 * clk_period;
	ASSERT (s_op1 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op2 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op3 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op4 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op5 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_final_output = 130) REPORT "the output should be '130'" SEVERITY ERROR;
	REPORT "_______________________";


	--emptying the pipeline
	REPORT "Finishing up and emptying the pipeline completely [a=0,b=0,c=0,d=0,e=0]";
	s_a <= 0;
	s_b <= 0;
	s_c <= 0;
	s_d <= 0;
	s_e <= 0;
	WAIT FOR 1 * clk_period;
	ASSERT (s_op1 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op2 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op3 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op4 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_op5 = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	ASSERT (s_final_output = 0) REPORT "the output should be '0'" SEVERITY ERROR;
	REPORT "_______________________";

	WAIT;

END PROCESS stim_process;
END;
